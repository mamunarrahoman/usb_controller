
`timescale 1ns/1ps
module usb_controller_tb;

reg clk;
reg reset;
reg mode;
reg L;
reg R;
reg U;
reg D;
reg A;
reg B;
reg X;
reg Y;

wire  out_cordinate_S;
wire  out_operation_S;
wire  [7:0]out_cordinate_P;
wire  [3:0]out_operation_P;

usb_controller duf(clk,reset,mode,L,R,U,D,A,B,X,Y,out_cordinate_P,out_operation_P,out_cordinate_S,out_operation_S);

initial
begin
	clk=1'b0;
	forever #0.25 clk=~clk;
end
initial
begin
	#0 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0;
	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0;

//mode_0_parallel data communication(gamming mode)
	#2 reset=1'b0;mode=1'b0;L=1'b1;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Left(L)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b1;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Right(R)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b0;U=1'b1;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Up(U)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b1;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Down(D)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
		
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //break

	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b1;B=1'b0;X=1'b0;Y=1'b0; //Enter(A)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b1;X=1'b0;Y=1'b0; //Back(B)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b1;Y=1'b0; //Option(X)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b1; //Properties(Y)
	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset

	#2 reset=1'b1;mode=1'b0;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //break

//mode_1_Serial data communication(Navigation Mode)
	#2 reset=1'b0;mode=1'b1;L=1'b1;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Left(L)
	#4
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b1;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Right(R)
	#4
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b0;U=1'b1;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Up(U)
	#3.75
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b1;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //Down(D)
	#6.25
	
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b0;U=1'b1;D=1'b1;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //marginal state check	
	
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset

	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //break

	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b1;B=1'b0;X=1'b0;Y=1'b0; //Enter(A)
	#4.75
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b1;X=1'b0;Y=1'b0; //Back(B)
	#5
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b1;Y=1'b0; //Option(X)
	#5
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	#2 reset=1'b0;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b1; //Properties(Y)
	#5
	#2 reset=1'b1;mode=1'b1;L=1'b0;R=1'b0;U=1'b0;D=1'b0;A=1'b0;B=1'b0;X=1'b0;Y=1'b0; //reset
	
	$finish;	

end
endmodule
